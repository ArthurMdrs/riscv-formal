// NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE
// This is an automatically generated file by arthur_linux on Wed Feb 21 13:03:42 -03 2024
//
// cmd:    veer -target=default -set build_axi4 
//

`include "common_defines.vh"
`undef TEC_RV_ICG
`define RV_PHYSICAL 1
